module top(
	input 			sys_clk,
	input 			rst_n,

	// 视频源输入
	// input 			video_clk, 
	// input 			video_rst, 
	// input 			video_de, 
	// input 	[15:0]	video_data0, 
	// input 	[15:0]	video_data1, 

	// 串口监测端口
	output 			uart_tx,
	output reg [23:0] rd_cnt,wr_cnt,

	// GMII输出
	output 			GMII_RST_N,
	output 			GMII_GTXCLK,
	output 			GMII_TXEN,
	output 			GMII_TXER,
	output 	[7:0]	GMII_TXD
	);

//此处使用RGB模拟一个1080P@30的时序
wire video_clk;
video_pll video_pll_m0(
	.clkin 	(sys_clk 		),
	.clkout (video_clk 		)
);

wire			video_rst; 
wire			video_de; 
wire	[15:0]	video_data; 
rgb1080P_sim rgb1080P_sim_m0(
	.sys_clk 			(video_clk 			),
	.rst_n 				(rst_n 				),

	.video_clk 			(video_clk 			),
	.video_de 			(video_de 			),
	.video_rst 			(video_rst 			),
	.video_data 		(video_data 		)
);

/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//////////////////// 			      接收模块	      	   /////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
wire [ 7:0] video_rd_data;
wire 		video_rd_en;

video_recive video_recive_m0(
	.Reset  			(video_rst			),
	
	.video_clk 			(video_clk 			),
	.video_de 			(video_de 			),
	.video_data 		(video_data 		),

	.video_rd_clk 		(GMII_GTXCLK 		),
	.video_rd_rdy 		(video_rd_rdy 		),
	.video_rd_en 		(video_rd_en 		),
	.video_rd_data 		(video_rd_data 		)
	);

/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//////////////////// 			      压缩模块	      	   /////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//未使用

/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//////////////////// 			      发送模块	      	   /////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
parameter DATA_SIZE = 16'D1442; // 2字节编号 + 1440字节数据
assign GMII_RST_N = rst_n;

GMII_pll GMII_pll_m0(
	.clkin 		(sys_clk 		), 
	.clkout  	(GMII_GTXCLK 	) // 125MHz
	);

wire send_start;
assign send_start   	= video_rd_rdy; // video_rd_num >= 1440;//(DATA_SIZE - 2); //当存满的数据足够一次发送，就开始发送(-2 编号字节) 
GMII_send #(
	.BOARD_MAC 	(48'h00_11_22_33_44_55 			),//开发板MAC地址
	.BOARD_IP 	({8'd192,8'd168,8'd1,8'd123}	),//开发板IP地址
	.BOARD_PORT (16'd8000 						),
	.DES_MAC 	(48'hff_ff_ff_ff_ff_ff 			),//目的MAC地址
	.DES_IP 	({8'd192,8'd168,8'd1,8'd102} 	),//目的IP地址
	.DES_PORT 	(16'd8001 						), //DES_PORT 
	.DATA_SIZE	(DATA_SIZE 						) //数据包长度 50~1500 B
	)GMII_send_m0(
	.rst_n 				(rst_n 				),

	.sys_clk 			(sys_clk 			),
	.frame_rst 			(video_rst 			),

	.send_start 		(send_start 		),
	.fifo_send_req 		(video_rd_en 		), 		
	.fifo_send_data 	(video_rd_data 		), 		

	.GMII_GTXCLK 		(GMII_GTXCLK 		),
	.GMII_TXD 			(GMII_TXD 			),
	.GMII_TXEN 			(GMII_TXEN 			),
	.GMII_TXER 			(GMII_TXER 			)
	);
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//////////////////// 			      监测模块	      	   /////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
always@(posedge GMII_GTXCLK) rd_cnt <=(!rst_n | video_rst)? 0 : video_rd_en? rd_cnt + 1 :rd_cnt ;
always@(posedge video_clk) wr_cnt 	<=(!rst_n | video_rst)? 0 : video_de? wr_cnt + 1 :wr_cnt ;


endmodule